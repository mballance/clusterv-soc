/****************************************************************************
 * clusterv_periph_subsys.v
 ****************************************************************************/
`include "wishbone_macros.svh"
  
/**
 * Module: clusterv_periph_subsys
 * 
 * TODO: Add module documentation
 */
module clusterv_periph_subsys(
		input				clock,
		input				reset);


endmodule


