/****************************************************************************
 * clusterv_soc.v
 ****************************************************************************/

/**
 * Module: clusterv_soc
 * 
 * TODO: Add module documentation
 */
module clusterv_soc(
		input		clock,
		input		reset
		);


endmodule


